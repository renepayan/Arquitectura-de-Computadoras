module vinculo (D,Q);
	input [7:0] D;
	input [7:0] Q;
	
	assign Q = D;
endmodule
