module vinculo (D,Q);
	input [7:0]: D;
	